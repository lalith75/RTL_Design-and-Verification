module clock_buffer(out,x);
input x;
output out;
buf b1(out,x);
endmodule
